module ycc_col_conv_g (data_a, data_b, result);
input wire [31:0] data_a; // this is the y input
input wire [31:0] data_b; // this is the CR value
output wire [31:0] result;

reg signed [31:0] temp1;
reg signed [31:0] temp2;
reg signed [31:0] cbg_val [255:0];
reg signed [31:0] crg_val [255:0];

always @(*) begin
	temp1 = (cbg_val[data_b[15:8]] + crg_val[data_b[7:0]]); //Sign extended right shift
	temp2 = (temp1[31] == 1) ? data_a-(~temp1+1) : data_a + temp1; //Sign extended right shift
	result = temp1;
end

always @(*) begin
crg_val[0] <= 32'h005b6900;
cbg_val[0] <= 32'h002c8d00;
crg_val[1] <= 32'h005ab22e;
cbg_val[1] <= 32'h002c34e6;
crg_val[2] <= 32'h0059fb5c;
cbg_val[2] <= 32'h002bdccc;
crg_val[3] <= 32'h0059448a;
cbg_val[3] <= 32'h002b84b2;
crg_val[4] <= 32'h00588db8;
cbg_val[4] <= 32'h002b2c98;
crg_val[5] <= 32'h0057d6e6;
cbg_val[5] <= 32'h002ad47e;
crg_val[6] <= 32'h00572014;
cbg_val[6] <= 32'h002a7c64;
crg_val[7] <= 32'h00566942;
cbg_val[7] <= 32'h002a244a;
crg_val[8] <= 32'h0055b270;
cbg_val[8] <= 32'h0029cc30;
crg_val[9] <= 32'h0054fb9e;
cbg_val[9] <= 32'h00297416;
crg_val[10] <= 32'h005444cc;
cbg_val[10] <= 32'h00291bfc;
crg_val[11] <= 32'h00538dfa;
cbg_val[11] <= 32'h0028c3e2;
crg_val[12] <= 32'h0052d728;
cbg_val[12] <= 32'h00286bc8;
crg_val[13] <= 32'h00522056;
cbg_val[13] <= 32'h002813ae;
crg_val[14] <= 32'h00516984;
cbg_val[14] <= 32'h0027bb94;
crg_val[15] <= 32'h0050b2b2;
cbg_val[15] <= 32'h0027637a;
crg_val[16] <= 32'h004ffbe0;
cbg_val[16] <= 32'h00270b60;
crg_val[17] <= 32'h004f450e;
cbg_val[17] <= 32'h0026b346;
crg_val[18] <= 32'h004e8e3c;
cbg_val[18] <= 32'h00265b2c;
crg_val[19] <= 32'h004dd76a;
cbg_val[19] <= 32'h00260312;
crg_val[20] <= 32'h004d2098;
cbg_val[20] <= 32'h0025aaf8;
crg_val[21] <= 32'h004c69c6;
cbg_val[21] <= 32'h002552de;
crg_val[22] <= 32'h004bb2f4;
cbg_val[22] <= 32'h0024fac4;
crg_val[23] <= 32'h004afc22;
cbg_val[23] <= 32'h0024a2aa;
crg_val[24] <= 32'h004a4550;
cbg_val[24] <= 32'h00244a90;
crg_val[25] <= 32'h00498e7e;
cbg_val[25] <= 32'h0023f276;
crg_val[26] <= 32'h0048d7ac;
cbg_val[26] <= 32'h00239a5c;
crg_val[27] <= 32'h004820da;
cbg_val[27] <= 32'h00234242;
crg_val[28] <= 32'h00476a08;
cbg_val[28] <= 32'h0022ea28;
crg_val[29] <= 32'h0046b336;
cbg_val[29] <= 32'h0022920e;
crg_val[30] <= 32'h0045fc64;
cbg_val[30] <= 32'h002239f4;
crg_val[31] <= 32'h00454592;
cbg_val[31] <= 32'h0021e1da;
crg_val[32] <= 32'h00448ec0;
cbg_val[32] <= 32'h002189c0;
crg_val[33] <= 32'h0043d7ee;
cbg_val[33] <= 32'h002131a6;
crg_val[34] <= 32'h0043211c;
cbg_val[34] <= 32'h0020d98c;
crg_val[35] <= 32'h00426a4a;
cbg_val[35] <= 32'h00208172;
crg_val[36] <= 32'h0041b378;
cbg_val[36] <= 32'h00202958;
crg_val[37] <= 32'h0040fca6;
cbg_val[37] <= 32'h001fd13e;
crg_val[38] <= 32'h004045d4;
cbg_val[38] <= 32'h001f7924;
crg_val[39] <= 32'h003f8f02;
cbg_val[39] <= 32'h001f210a;
crg_val[40] <= 32'h003ed830;
cbg_val[40] <= 32'h001ec8f0;
crg_val[41] <= 32'h003e215e;
cbg_val[41] <= 32'h001e70d6;
crg_val[42] <= 32'h003d6a8c;
cbg_val[42] <= 32'h001e18bc;
crg_val[43] <= 32'h003cb3ba;
cbg_val[43] <= 32'h001dc0a2;
crg_val[44] <= 32'h003bfce8;
cbg_val[44] <= 32'h001d6888;
crg_val[45] <= 32'h003b4616;
cbg_val[45] <= 32'h001d106e;
crg_val[46] <= 32'h003a8f44;
cbg_val[46] <= 32'h001cb854;
crg_val[47] <= 32'h0039d872;
cbg_val[47] <= 32'h001c603a;
crg_val[48] <= 32'h003921a0;
cbg_val[48] <= 32'h001c0820;
crg_val[49] <= 32'h00386ace;
cbg_val[49] <= 32'h001bb006;
crg_val[50] <= 32'h0037b3fc;
cbg_val[50] <= 32'h001b57ec;
crg_val[51] <= 32'h0036fd2a;
cbg_val[51] <= 32'h001affd2;
crg_val[52] <= 32'h00364658;
cbg_val[52] <= 32'h001aa7b8;
crg_val[53] <= 32'h00358f86;
cbg_val[53] <= 32'h001a4f9e;
crg_val[54] <= 32'h0034d8b4;
cbg_val[54] <= 32'h0019f784;
crg_val[55] <= 32'h003421e2;
cbg_val[55] <= 32'h00199f6a;
crg_val[56] <= 32'h00336b10;
cbg_val[56] <= 32'h00194750;
crg_val[57] <= 32'h0032b43e;
cbg_val[57] <= 32'h0018ef36;
crg_val[58] <= 32'h0031fd6c;
cbg_val[58] <= 32'h0018971c;
crg_val[59] <= 32'h0031469a;
cbg_val[59] <= 32'h00183f02;
crg_val[60] <= 32'h00308fc8;
cbg_val[60] <= 32'h0017e6e8;
crg_val[61] <= 32'h002fd8f6;
cbg_val[61] <= 32'h00178ece;
crg_val[62] <= 32'h002f2224;
cbg_val[62] <= 32'h001736b4;
crg_val[63] <= 32'h002e6b52;
cbg_val[63] <= 32'h0016de9a;
crg_val[64] <= 32'h002db480;
cbg_val[64] <= 32'h00168680;
crg_val[65] <= 32'h002cfdae;
cbg_val[65] <= 32'h00162e66;
crg_val[66] <= 32'h002c46dc;
cbg_val[66] <= 32'h0015d64c;
crg_val[67] <= 32'h002b900a;
cbg_val[67] <= 32'h00157e32;
crg_val[68] <= 32'h002ad938;
cbg_val[68] <= 32'h00152618;
crg_val[69] <= 32'h002a2266;
cbg_val[69] <= 32'h0014cdfe;
crg_val[70] <= 32'h00296b94;
cbg_val[70] <= 32'h001475e4;
crg_val[71] <= 32'h0028b4c2;
cbg_val[71] <= 32'h00141dca;
crg_val[72] <= 32'h0027fdf0;
cbg_val[72] <= 32'h0013c5b0;
crg_val[73] <= 32'h0027471e;
cbg_val[73] <= 32'h00136d96;
crg_val[74] <= 32'h0026904c;
cbg_val[74] <= 32'h0013157c;
crg_val[75] <= 32'h0025d97a;
cbg_val[75] <= 32'h0012bd62;
crg_val[76] <= 32'h002522a8;
cbg_val[76] <= 32'h00126548;
crg_val[77] <= 32'h00246bd6;
cbg_val[77] <= 32'h00120d2e;
crg_val[78] <= 32'h0023b504;
cbg_val[78] <= 32'h0011b514;
crg_val[79] <= 32'h0022fe32;
cbg_val[79] <= 32'h00115cfa;
crg_val[80] <= 32'h00224760;
cbg_val[80] <= 32'h001104e0;
crg_val[81] <= 32'h0021908e;
cbg_val[81] <= 32'h0010acc6;
crg_val[82] <= 32'h0020d9bc;
cbg_val[82] <= 32'h001054ac;
crg_val[83] <= 32'h002022ea;
cbg_val[83] <= 32'h000ffc92;
crg_val[84] <= 32'h001f6c18;
cbg_val[84] <= 32'h000fa478;
crg_val[85] <= 32'h001eb546;
cbg_val[85] <= 32'h000f4c5e;
crg_val[86] <= 32'h001dfe74;
cbg_val[86] <= 32'h000ef444;
crg_val[87] <= 32'h001d47a2;
cbg_val[87] <= 32'h000e9c2a;
crg_val[88] <= 32'h001c90d0;
cbg_val[88] <= 32'h000e4410;
crg_val[89] <= 32'h001bd9fe;
cbg_val[89] <= 32'h000debf6;
crg_val[90] <= 32'h001b232c;
cbg_val[90] <= 32'h000d93dc;
crg_val[91] <= 32'h001a6c5a;
cbg_val[91] <= 32'h000d3bc2;
crg_val[92] <= 32'h0019b588;
cbg_val[92] <= 32'h000ce3a8;
crg_val[93] <= 32'h0018feb6;
cbg_val[93] <= 32'h000c8b8e;
crg_val[94] <= 32'h001847e4;
cbg_val[94] <= 32'h000c3374;
crg_val[95] <= 32'h00179112;
cbg_val[95] <= 32'h000bdb5a;
crg_val[96] <= 32'h0016da40;
cbg_val[96] <= 32'h000b8340;
crg_val[97] <= 32'h0016236e;
cbg_val[97] <= 32'h000b2b26;
crg_val[98] <= 32'h00156c9c;
cbg_val[98] <= 32'h000ad30c;
crg_val[99] <= 32'h0014b5ca;
cbg_val[99] <= 32'h000a7af2;
crg_val[100] <= 32'h0013fef8;
cbg_val[100] <= 32'h000a22d8;
crg_val[101] <= 32'h00134826;
cbg_val[101] <= 32'h0009cabe;
crg_val[102] <= 32'h00129154;
cbg_val[102] <= 32'h000972a4;
crg_val[103] <= 32'h0011da82;
cbg_val[103] <= 32'h00091a8a;
crg_val[104] <= 32'h001123b0;
cbg_val[104] <= 32'h0008c270;
crg_val[105] <= 32'h00106cde;
cbg_val[105] <= 32'h00086a56;
crg_val[106] <= 32'h000fb60c;
cbg_val[106] <= 32'h0008123c;
crg_val[107] <= 32'h000eff3a;
cbg_val[107] <= 32'h0007ba22;
crg_val[108] <= 32'h000e4868;
cbg_val[108] <= 32'h00076208;
crg_val[109] <= 32'h000d9196;
cbg_val[109] <= 32'h000709ee;
crg_val[110] <= 32'h000cdac4;
cbg_val[110] <= 32'h0006b1d4;
crg_val[111] <= 32'h000c23f2;
cbg_val[111] <= 32'h000659ba;
crg_val[112] <= 32'h000b6d20;
cbg_val[112] <= 32'h000601a0;
crg_val[113] <= 32'h000ab64e;
cbg_val[113] <= 32'h0005a986;
crg_val[114] <= 32'h0009ff7c;
cbg_val[114] <= 32'h0005516c;
crg_val[115] <= 32'h000948aa;
cbg_val[115] <= 32'h0004f952;
crg_val[116] <= 32'h000891d8;
cbg_val[116] <= 32'h0004a138;
crg_val[117] <= 32'h0007db06;
cbg_val[117] <= 32'h0004491e;
crg_val[118] <= 32'h00072434;
cbg_val[118] <= 32'h0003f104;
crg_val[119] <= 32'h00066d62;
cbg_val[119] <= 32'h000398ea;
crg_val[120] <= 32'h0005b690;
cbg_val[120] <= 32'h000340d0;
crg_val[121] <= 32'h0004ffbe;
cbg_val[121] <= 32'h0002e8b6;
crg_val[122] <= 32'h000448ec;
cbg_val[122] <= 32'h0002909c;
crg_val[123] <= 32'h0003921a;
cbg_val[123] <= 32'h00023882;
crg_val[124] <= 32'h0002db48;
cbg_val[124] <= 32'h0001e068;
crg_val[125] <= 32'h00022476;
cbg_val[125] <= 32'h0001884e;
crg_val[126] <= 32'h00016da4;
cbg_val[126] <= 32'h00013034;
crg_val[127] <= 32'h0000b6d2;
cbg_val[127] <= 32'h0000d81a;
crg_val[128] <= 32'h00000000;
cbg_val[128] <= 32'h00008000;
crg_val[129] <= 32'hffff492e;
cbg_val[129] <= 32'h000027e6;
crg_val[130] <= 32'hfffe925c;
cbg_val[130] <= 32'hffffcfcc;
crg_val[131] <= 32'hfffddb8a;
cbg_val[131] <= 32'hffff77b2;
crg_val[132] <= 32'hfffd24b8;
cbg_val[132] <= 32'hffff1f98;
crg_val[133] <= 32'hfffc6de6;
cbg_val[133] <= 32'hfffec77e;
crg_val[134] <= 32'hfffbb714;
cbg_val[134] <= 32'hfffe6f64;
crg_val[135] <= 32'hfffb0042;
cbg_val[135] <= 32'hfffe174a;
crg_val[136] <= 32'hfffa4970;
cbg_val[136] <= 32'hfffdbf30;
crg_val[137] <= 32'hfff9929e;
cbg_val[137] <= 32'hfffd6716;
crg_val[138] <= 32'hfff8dbcc;
cbg_val[138] <= 32'hfffd0efc;
crg_val[139] <= 32'hfff824fa;
cbg_val[139] <= 32'hfffcb6e2;
crg_val[140] <= 32'hfff76e28;
cbg_val[140] <= 32'hfffc5ec8;
crg_val[141] <= 32'hfff6b756;
cbg_val[141] <= 32'hfffc06ae;
crg_val[142] <= 32'hfff60084;
cbg_val[142] <= 32'hfffbae94;
crg_val[143] <= 32'hfff549b2;
cbg_val[143] <= 32'hfffb567a;
crg_val[144] <= 32'hfff492e0;
cbg_val[144] <= 32'hfffafe60;
crg_val[145] <= 32'hfff3dc0e;
cbg_val[145] <= 32'hfffaa646;
crg_val[146] <= 32'hfff3253c;
cbg_val[146] <= 32'hfffa4e2c;
crg_val[147] <= 32'hfff26e6a;
cbg_val[147] <= 32'hfff9f612;
crg_val[148] <= 32'hfff1b798;
cbg_val[148] <= 32'hfff99df8;
crg_val[149] <= 32'hfff100c6;
cbg_val[149] <= 32'hfff945de;
crg_val[150] <= 32'hfff049f4;
cbg_val[150] <= 32'hfff8edc4;
crg_val[151] <= 32'hffef9322;
cbg_val[151] <= 32'hfff895aa;
crg_val[152] <= 32'hffeedc50;
cbg_val[152] <= 32'hfff83d90;
crg_val[153] <= 32'hffee257e;
cbg_val[153] <= 32'hfff7e576;
crg_val[154] <= 32'hffed6eac;
cbg_val[154] <= 32'hfff78d5c;
crg_val[155] <= 32'hffecb7da;
cbg_val[155] <= 32'hfff73542;
crg_val[156] <= 32'hffec0108;
cbg_val[156] <= 32'hfff6dd28;
crg_val[157] <= 32'hffeb4a36;
cbg_val[157] <= 32'hfff6850e;
crg_val[158] <= 32'hffea9364;
cbg_val[158] <= 32'hfff62cf4;
crg_val[159] <= 32'hffe9dc92;
cbg_val[159] <= 32'hfff5d4da;
crg_val[160] <= 32'hffe925c0;
cbg_val[160] <= 32'hfff57cc0;
crg_val[161] <= 32'hffe86eee;
cbg_val[161] <= 32'hfff524a6;
crg_val[162] <= 32'hffe7b81c;
cbg_val[162] <= 32'hfff4cc8c;
crg_val[163] <= 32'hffe7014a;
cbg_val[163] <= 32'hfff47472;
crg_val[164] <= 32'hffe64a78;
cbg_val[164] <= 32'hfff41c58;
crg_val[165] <= 32'hffe593a6;
cbg_val[165] <= 32'hfff3c43e;
crg_val[166] <= 32'hffe4dcd4;
cbg_val[166] <= 32'hfff36c24;
crg_val[167] <= 32'hffe42602;
cbg_val[167] <= 32'hfff3140a;
crg_val[168] <= 32'hffe36f30;
cbg_val[168] <= 32'hfff2bbf0;
crg_val[169] <= 32'hffe2b85e;
cbg_val[169] <= 32'hfff263d6;
crg_val[170] <= 32'hffe2018c;
cbg_val[170] <= 32'hfff20bbc;
crg_val[171] <= 32'hffe14aba;
cbg_val[171] <= 32'hfff1b3a2;
crg_val[172] <= 32'hffe093e8;
cbg_val[172] <= 32'hfff15b88;
crg_val[173] <= 32'hffdfdd16;
cbg_val[173] <= 32'hfff1036e;
crg_val[174] <= 32'hffdf2644;
cbg_val[174] <= 32'hfff0ab54;
crg_val[175] <= 32'hffde6f72;
cbg_val[175] <= 32'hfff0533a;
crg_val[176] <= 32'hffddb8a0;
cbg_val[176] <= 32'hffeffb20;
crg_val[177] <= 32'hffdd01ce;
cbg_val[177] <= 32'hffefa306;
crg_val[178] <= 32'hffdc4afc;
cbg_val[178] <= 32'hffef4aec;
crg_val[179] <= 32'hffdb942a;
cbg_val[179] <= 32'hffeef2d2;
crg_val[180] <= 32'hffdadd58;
cbg_val[180] <= 32'hffee9ab8;
crg_val[181] <= 32'hffda2686;
cbg_val[181] <= 32'hffee429e;
crg_val[182] <= 32'hffd96fb4;
cbg_val[182] <= 32'hffedea84;
crg_val[183] <= 32'hffd8b8e2;
cbg_val[183] <= 32'hffed926a;
crg_val[184] <= 32'hffd80210;
cbg_val[184] <= 32'hffed3a50;
crg_val[185] <= 32'hffd74b3e;
cbg_val[185] <= 32'hffece236;
crg_val[186] <= 32'hffd6946c;
cbg_val[186] <= 32'hffec8a1c;
crg_val[187] <= 32'hffd5dd9a;
cbg_val[187] <= 32'hffec3202;
crg_val[188] <= 32'hffd526c8;
cbg_val[188] <= 32'hffebd9e8;
crg_val[189] <= 32'hffd46ff6;
cbg_val[189] <= 32'hffeb81ce;
crg_val[190] <= 32'hffd3b924;
cbg_val[190] <= 32'hffeb29b4;
crg_val[191] <= 32'hffd30252;
cbg_val[191] <= 32'hffead19a;
crg_val[192] <= 32'hffd24b80;
cbg_val[192] <= 32'hffea7980;
crg_val[193] <= 32'hffd194ae;
cbg_val[193] <= 32'hffea2166;
crg_val[194] <= 32'hffd0dddc;
cbg_val[194] <= 32'hffe9c94c;
crg_val[195] <= 32'hffd0270a;
cbg_val[195] <= 32'hffe97132;
crg_val[196] <= 32'hffcf7038;
cbg_val[196] <= 32'hffe91918;
crg_val[197] <= 32'hffceb966;
cbg_val[197] <= 32'hffe8c0fe;
crg_val[198] <= 32'hffce0294;
cbg_val[198] <= 32'hffe868e4;
crg_val[199] <= 32'hffcd4bc2;
cbg_val[199] <= 32'hffe810ca;
crg_val[200] <= 32'hffcc94f0;
cbg_val[200] <= 32'hffe7b8b0;
crg_val[201] <= 32'hffcbde1e;
cbg_val[201] <= 32'hffe76096;
crg_val[202] <= 32'hffcb274c;
cbg_val[202] <= 32'hffe7087c;
crg_val[203] <= 32'hffca707a;
cbg_val[203] <= 32'hffe6b062;
crg_val[204] <= 32'hffc9b9a8;
cbg_val[204] <= 32'hffe65848;
crg_val[205] <= 32'hffc902d6;
cbg_val[205] <= 32'hffe6002e;
crg_val[206] <= 32'hffc84c04;
cbg_val[206] <= 32'hffe5a814;
crg_val[207] <= 32'hffc79532;
cbg_val[207] <= 32'hffe54ffa;
crg_val[208] <= 32'hffc6de60;
cbg_val[208] <= 32'hffe4f7e0;
crg_val[209] <= 32'hffc6278e;
cbg_val[209] <= 32'hffe49fc6;
crg_val[210] <= 32'hffc570bc;
cbg_val[210] <= 32'hffe447ac;
crg_val[211] <= 32'hffc4b9ea;
cbg_val[211] <= 32'hffe3ef92;
crg_val[212] <= 32'hffc40318;
cbg_val[212] <= 32'hffe39778;
crg_val[213] <= 32'hffc34c46;
cbg_val[213] <= 32'hffe33f5e;
crg_val[214] <= 32'hffc29574;
cbg_val[214] <= 32'hffe2e744;
crg_val[215] <= 32'hffc1dea2;
cbg_val[215] <= 32'hffe28f2a;
crg_val[216] <= 32'hffc127d0;
cbg_val[216] <= 32'hffe23710;
crg_val[217] <= 32'hffc070fe;
cbg_val[217] <= 32'hffe1def6;
crg_val[218] <= 32'hffbfba2c;
cbg_val[218] <= 32'hffe186dc;
crg_val[219] <= 32'hffbf035a;
cbg_val[219] <= 32'hffe12ec2;
crg_val[220] <= 32'hffbe4c88;
cbg_val[220] <= 32'hffe0d6a8;
crg_val[221] <= 32'hffbd95b6;
cbg_val[221] <= 32'hffe07e8e;
crg_val[222] <= 32'hffbcdee4;
cbg_val[222] <= 32'hffe02674;
crg_val[223] <= 32'hffbc2812;
cbg_val[223] <= 32'hffdfce5a;
crg_val[224] <= 32'hffbb7140;
cbg_val[224] <= 32'hffdf7640;
crg_val[225] <= 32'hffbaba6e;
cbg_val[225] <= 32'hffdf1e26;
crg_val[226] <= 32'hffba039c;
cbg_val[226] <= 32'hffdec60c;
crg_val[227] <= 32'hffb94cca;
cbg_val[227] <= 32'hffde6df2;
crg_val[228] <= 32'hffb895f8;
cbg_val[228] <= 32'hffde15d8;
crg_val[229] <= 32'hffb7df26;
cbg_val[229] <= 32'hffddbdbe;
crg_val[230] <= 32'hffb72854;
cbg_val[230] <= 32'hffdd65a4;
crg_val[231] <= 32'hffb67182;
cbg_val[231] <= 32'hffdd0d8a;
crg_val[232] <= 32'hffb5bab0;
cbg_val[232] <= 32'hffdcb570;
crg_val[233] <= 32'hffb503de;
cbg_val[233] <= 32'hffdc5d56;
crg_val[234] <= 32'hffb44d0c;
cbg_val[234] <= 32'hffdc053c;
crg_val[235] <= 32'hffb3963a;
cbg_val[235] <= 32'hffdbad22;
crg_val[236] <= 32'hffb2df68;
cbg_val[236] <= 32'hffdb5508;
crg_val[237] <= 32'hffb22896;
cbg_val[237] <= 32'hffdafcee;
crg_val[238] <= 32'hffb171c4;
cbg_val[238] <= 32'hffdaa4d4;
crg_val[239] <= 32'hffb0baf2;
cbg_val[239] <= 32'hffda4cba;
crg_val[240] <= 32'hffb00420;
cbg_val[240] <= 32'hffd9f4a0;
crg_val[241] <= 32'hffaf4d4e;
cbg_val[241] <= 32'hffd99c86;
crg_val[242] <= 32'hffae967c;
cbg_val[242] <= 32'hffd9446c;
crg_val[243] <= 32'hffaddfaa;
cbg_val[243] <= 32'hffd8ec52;
crg_val[244] <= 32'hffad28d8;
cbg_val[244] <= 32'hffd89438;
crg_val[245] <= 32'hffac7206;
cbg_val[245] <= 32'hffd83c1e;
crg_val[246] <= 32'hffabbb34;
cbg_val[246] <= 32'hffd7e404;
crg_val[247] <= 32'hffab0462;
cbg_val[247] <= 32'hffd78bea;
crg_val[248] <= 32'hffaa4d90;
cbg_val[248] <= 32'hffd733d0;
crg_val[249] <= 32'hffa996be;
cbg_val[249] <= 32'hffd6dbb6;
crg_val[250] <= 32'hffa8dfec;
cbg_val[250] <= 32'hffd6839c;
crg_val[251] <= 32'hffa8291a;
cbg_val[251] <= 32'hffd62b82;
crg_val[252] <= 32'hffa77248;
cbg_val[252] <= 32'hffd5d368;
crg_val[253] <= 32'hffa6bb76;
cbg_val[253] <= 32'hffd57b4e;
crg_val[254] <= 32'hffa604a4;
cbg_val[254] <= 32'hffd52334;
crg_val[255] <= 32'hffa54dd2;
cbg_val[255] <= 32'hffd4cb1a;
end

endmodule
